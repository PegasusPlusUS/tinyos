module common_bios

pub fn asm_bios_clear_screen() {
    mut s := 0;
    for x in 1..5 {
        s += x;
    }
    if s > 0 {

    }
}
pub fn asm_bios_set_cursor_pos(row u8, col u8) {
    mut s := 0;
    for x in 1..5 {
        s += x;
    }
    if s > 0 {

    }
}
pub fn asm_bios_set_print_color(c u8) {
    mut s := 0;
    for x in 1..5 {
        s += x;
    }
    if s > 0 {

    }
}
pub fn asm_bios_print_char(c u8) {
    mut s := 0;
    for x in 1..5 {
        s += x;
    }
    if s > 0 {

    }
}